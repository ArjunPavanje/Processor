`include "shift/shift.v"
`include "addsub/addsub.v"
`include "mul/mul.v"

module FPMul (
    input  [63:0] N1,
    input  [63:0] N2,
    output [63:0] out
);

  // Extracting Sign, Exponent, Mantissa
  wire [51:0] M_1;
  wire [51:0] M_2;
  wire [10:0] E_1;
  wire [10:0] E_2;
  wire S_1;
  wire S_2;
  assign M_1 = N1[51:0];
  assign M_2 = N2[51:0];

  assign E_1 = N1[62:52];
  assign E_2 = N2[62:52];

  assign S_1 = N1[63];
  assign S_2 = N2[63];


  wire [63:0] temp1;
  wire [63:0] temp2;
  assign temp1 = {12'b1, M_1};
  assign temp2 = {12'b1, M_2};
  // Multiplying mantissas M_1 and M_2
  wire [127:0] mantissa_product;
  mul FPmul_mantissa (
      .a({12'b1, M_1}),
      .b({12'b1, M_2}),
      .sign(1'b0),
      .res(mantissa_product)
  );
  // Normalizing mantissa
  wire [52:0] mantissa_normalized;
  wire L;
  wire G;
  wire R;
  wire S;
  wire round;

  // Also setting LSB, Guard, Round, Sticky bits
  assign mantissa_normalized = (mantissa_product[105])?mantissa_product[105:53]:mantissa_product[104:52];
  assign L = (mantissa_product[105]) ? mantissa_product[53] : mantissa_product[52];
  assign G = (mantissa_product[105]) ? mantissa_product[52] : mantissa_product[51];
  assign R = (mantissa_product[105]) ? mantissa_product[51] : mantissa_product[50];
  assign S = (mantissa_product[105]) ? |mantissa_product[50:0] : |mantissa_product[49:0];

  assign round = (G & (R | S)) | (L & G & (~R) & (~S));

  wire [63:0] mantissa_rounded;
  wire cout;
  addsub FPmul_round (
      .a({11'b0, mantissa_normalized}),
      .b((round) ? {63'b0, 1'b1} : {63'b0, 1'b0}),
      .sel(1'b0),
      .cout(cout),
      .res(mantissa_rounded)
  );

  wire [51:0] mantissa_renormalized;
  assign mantissa_renormalized = (cout) ? mantissa_rounded[52:1] : mantissa_rounded[51:0];
  assign out[51:0] = mantissa_renormalized;
  assign out[63:52] = 12'b0;

endmodule
